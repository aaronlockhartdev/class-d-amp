.SUBCKT Lead_14 1 2
R1 7 1 1
C1 6 1 1
C2 7 6 1
C3 2 3 1
C4 3 7 1
R2 2 7 1
R3 0 6 1
R4 0 7 1
R5 0 3 1
.ENDS
