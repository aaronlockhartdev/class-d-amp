C:\Users\Aaron\Documents\GitHub\class-d-amp\loop_analysis\sym_analysis\SapWin\class_d_4.sch
R1 1 0 1
R2 7 1 1
EO1 3 0 1 0 1e6
C1 3 1 1
C2 4 2 1
EO2 4 0 2 0 1e6
R3 2 3 1
R4 10 4 1
V1 5 0 AC 1
L1 7 5 1
C4 7 0 1
R7 7 0 4
R10 6 11 1
C7 6 7 1
R9 0 8 1
C6 8 7 1
R8 0 9 1
C5 8 9 1
C3 9 11 1
R6 10 11 1
.AC DEC 100 1 1000
.PROBE
.END
