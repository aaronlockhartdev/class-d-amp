C:\Users\Aaron\Documents\GitHub\class-d-amp\SapWin\Class-D MFB.sch
Rg1 7 1 1
Ri 1 0 1800
Rfb 1 5 8200
EO2 0 0 7 0 1e6
Cmfb1 9 0 1e-10
Rmfb 3 2 680
EO1 2 0 8 0 1e6
Cmfb2 2 8 1e-09
Rmfb3 2 9 2200
Rload 5 0 4
Rl 4 5 1000
Cl 3 4 3.3e-10
Cf 5 0 6.8e-07
Lf 5 6 1e-05
V1 6 0 AC 1
Rg2 0 7 1
Rmfb2 8 9 1
Rmfb1 9 0 1
.AC DEC 100 1 1000
.PROBE
.END
