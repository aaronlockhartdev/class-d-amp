.SUBCKT MFB 1 2
R1 5 1 1
R2 6 5 1
C1 0 5 1
C2 6 2 1
R1 5 2 1
EO1 2 0 6 0 1e6
.ENDS
